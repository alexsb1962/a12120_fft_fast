library verilog;
use verilog.vl_types.all;
entity fast_fft_tb is
end fast_fft_tb;

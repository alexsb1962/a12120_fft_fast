library verilog;
use verilog.vl_types.all;
entity dsp_tb is
end dsp_tb;

library verilog;
use verilog.vl_types.all;
entity fifo_120_48_tb is
end fifo_120_48_tb;
